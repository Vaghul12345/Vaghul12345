module datapath(clk, Alu,
